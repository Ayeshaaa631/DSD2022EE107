module segment(
    input a1,a0,b1,b0,x,y,z,
    output reg SegA, SegB, SegC, SegD, SegE, SegF, SegG, An0, An1, An2, An3, An4, An5, An6, An7
);
always @(*) begin
    An0 = ((x)||(y)||(z));
    An1 = ((x)||(y)||(~z));
    An2 = ((x)||(~y)||(z));
    An3 = ((x)||(~y)||(~z));
    An4 = ((~x)||(y)||(z));
    An5 = ((~x)||(y)||(~z));
    An6 = ((~x)||(~y)||(z));
    An7 = ((~x)||(~y)||(~z));
    SegA = ((~a1)&&(~a0)&&(~b1)&&(b0))||((~a1)&&(a0)&&(~b1)&&(~b0))||((a1)&&(a0)&&(~b1)&&(b0))||((a1)&&(~a0)&&(b1)&&(b0));
    SegB = ((a1)&&(b1)&&(b0))||((a0)&&(b1)&&(~b0))||((a1)&&(a0)&&(~b0))||((~a1)&&(a0)&&(~b1)&&(b0));
    SegC = ((a1)&&(a0)&&(~b0))||((a1)&&(a0)&&(b1))||((~a1)&&(~a0)&&(b1)&&(~b0));
    SegD = ((a0)&&(b1)&&(b0))||((~a1)&&(a0)&&(~b1)&&(~b0))||((~a1)&&(~a0)&&(~b1)&&(b0))||((a1)&&(~a0)&&(b1)&&(~b0));
    SegE = ((~a1)&&(a0)&&(~b1))||((~a1)&&(b0))||((~a0)&&(~b1)&&(b0));
    SegF = ((~a1)&&(b1)&&(b0))||((~a1)&&(~a0)&&(b0))||((~a1)&&(~a0)&&(b1))||((a1)&&(a0)&&(~b1)&&(b0));
    SegG = ((~a1)&&(~a0)&&(~b1))||((a1)&&(a0)&&(~b1)&&(~b0))||((~a1)&&(a0)&&(b1)&&(b0));
end
endmodule
